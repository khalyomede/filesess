module filesess

pub struct SessionData {
	value string
	flashed bool
}
